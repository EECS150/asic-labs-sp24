`include "alu_op.vh"

module alu(
    input [31:0] a, b,
    input [3:0] alu_op,
    output [31:0] out
);

// Your code goes here

endmodule
